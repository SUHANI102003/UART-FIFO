`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 01.09.2024 10:51:38
// Design Name: 
// Module Name: debouncer_delayed_fsm
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module debouncer_delayed_fsm(
 input clk,reset_n,
 input noisy,timer_done,
 output debounce, timer_reset
    );
 
 reg [1:0] state_next, state_reg;   
parameter s0 = 0, s1 = 1,  s2 = 2,  s3 = 3 ;
 
// state register
always@(posedge clk, negedge reset_n)
begin
    if(~reset_n)
        state_reg <= 0;
    else 
        state_reg <= state_next;
end

// next state logic
always@(*)
begin
    state_next = state_reg;
    case(state_reg)
    s0 : if(~noisy)
            state_next = s0;
         else
             state_next = s1;
    s1 : if(~noisy)
            state_next = s0;
         else if(noisy & ~timer_done)
             state_next = s1;
         else if(noisy & timer_done)
             state_next = s2;
    s2 : if(noisy)
            state_next = s2;
         else
             state_next = s3;
    s3 : if(noisy)
            state_next = s2;
         else if(~noisy & ~timer_done)
             state_next = s3;
         else if(~noisy & timer_done)
             state_next = s0;
    default : state_next = s0;
    
    endcase
end

//output logic
assign timer_reset = (state_reg == s0) | (state_reg == s2);
assign debounce = (state_reg == s2) | (state_reg == s3);
  
endmodule


/* This fsm code is designed in such a way that we need to 
set the timer according to the value we need.
So, what we can do is create a timer module and 
instantiate it in debounce fsm code

timer module is just a counter that ticks when 
value specified as time is reached
*/